** sch_path: /foss/designs/Assignment2/src/CS_Current_Mirror.sch
**.subckt CS_Current_Mirror vin vout vdd iref
*.ipin vin
*.opin vout
*.iopin vdd
*.iopin iref
XC1 vout GND sky130_fd_pr__cap_mim_m3_1 W=40 L=87 MF=1 m=1
XM2 vout iref vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=170 nf=15 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 vout vin GND GND sky130_fd_pr__nfet_01v8 L=1 W=120 nf=12 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 iref iref vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=170 nf=15 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt




.option temp=27
.option gmin = 1e-12
.param vbias = 0.7180

vdd vdd 0 1.8
*vin vin 0 dc {vbias} ac 0.1
vin vin 0 dc {vbias} ac 0.01 0 SIN({vbias} 0.01 100k)
iref iref 0 dc 0.327m

.dc vin 0 1.8 10m
.ac dec 10 10 200Meg


.tran 0.1u 20u 1n

.saveall
.control
run

setplot dc1
plot v(vin) v(vout) 0.9
plot -i(vdd) vs v(vin)


setplot ac1
plot db(v(vout)/v(vin))
*plot mag(ac1.v(vout))

setplot tran1
plot v(vin) v(vout)

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
